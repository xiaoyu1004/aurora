`ifndef GLOBAL_CONFIG_VH
`define GLOBAL_CONFIG_VH

`define ENABLE      1
`define DISABLE     0

`endif